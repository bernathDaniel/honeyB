//=============================================================================
// Project  : HoneyB V7
// File Name: top_seq_lib.sv
//=============================================================================
// Description: Sequence for top
// IMPORANT   : Right now the child sequences
//              are within a fork...join however
//              this might be changed to fork...join_none
//              In the case we might want multiple read/write operations.
//=============================================================================

`ifndef TOP_SEQ_LIB_SV
`define TOP_SEQ_LIB_SV

`include "uvm_macros.svh"
import uvm_pkg::*;
import honeyb_pkg::*;

class top_default_seq extends uvm_sequence #(uvm_sequence_item);

  `uvm_object_utils(top_default_seq)

  xlr_mem_agent  m_xlr_mem_agent;
  xlr_gpp_agent  m_xlr_gpp_agent;

  // Sequence #
  int m_seq_count = 5;

  // Sequence iteration counter
  int iteration_count = 0;

  extern function new(string name = "");
  extern task body();
  extern task pre_start();
  extern task post_start();

`ifndef UVM_POST_VERSION_1_1
  // Functions to support UVM 1.2 objection API in UVM 1.1
  extern function uvm_phase get_starting_phase();
  extern function void set_starting_phase(uvm_phase phase);
`endif

endclass : top_default_seq


function top_default_seq::new(string name = "");
  super.new(name);
endfunction : new


task top_default_seq::body();
  `honeyb("TOP SEQ", "New sequence starting...")

  repeat (m_seq_count)
  begin
    fork
      if (( m_xlr_mem_agent.m_config.is_active   == UVM_ACTIVE) &&
            m_xlr_mem_agent.m_config.mem_is_used == 1'b0            )
      begin
        xlr_mem_default_seq seq;
        seq = xlr_mem_default_seq::type_id::create("seq");
        seq.set_item_context(this, m_xlr_mem_agent.m_sequencer);
        if ( !seq.randomize() )
          `uvm_error("", "Failed to randomize sequence")
        seq.set_starting_phase( get_starting_phase() );
        seq.start(m_xlr_mem_agent.m_sequencer, this);        
      end else `honeyb("TOP SEQ", "MEM SEQ UNINITIALIZED ", "STATUS = OK")

      if (m_xlr_gpp_agent.m_config.is_active == UVM_ACTIVE)
      begin
        xlr_gpp_default_seq seq;
        seq = xlr_gpp_default_seq::type_id::create("seq");
        seq.set_item_context(this, m_xlr_gpp_agent.m_sequencer);
        if ( !seq.randomize() )
          `uvm_error("", "Failed to randomize sequence")
        seq.set_starting_phase( get_starting_phase() );
        seq.start(m_xlr_gpp_agent.m_sequencer, this);
      end
    join
  end

  `honeyb("TOP SEQ", "Sequence completed...")
endtask : body


task top_default_seq::pre_start();
  uvm_phase phase = get_starting_phase();
  if (phase != null)
    phase.raise_objection(this);
endtask: pre_start


task top_default_seq::post_start();
  uvm_phase phase = get_starting_phase();
  if (phase != null) 
    phase.drop_objection(this);
endtask: post_start


`ifndef UVM_POST_VERSION_1_1
  function uvm_phase top_default_seq::get_starting_phase();
    return starting_phase;
  endfunction: get_starting_phase


  function void top_default_seq::set_starting_phase(uvm_phase phase);
    starting_phase = phase;
  endfunction: set_starting_phase
`endif

`endif // TOP_SEQ_LIB_SV